library verilog;
use verilog.vl_types.all;
entity TDC_result is
    port(
        TDC_value_31    : out    vl_logic;
        TDC_value_30    : out    vl_logic;
        TDC_value_29    : out    vl_logic;
        TDC_value_28    : out    vl_logic;
        TDC_value_27    : out    vl_logic;
        TDC_value_26    : out    vl_logic;
        TDC_value_25    : out    vl_logic;
        TDC_value_24    : out    vl_logic;
        TDC_value_23    : out    vl_logic;
        TDC_value_22    : out    vl_logic;
        TDC_value_21    : out    vl_logic;
        TDC_value_20    : out    vl_logic;
        TDC_value_19    : out    vl_logic;
        TDC_value_18    : out    vl_logic;
        TDC_value_17    : out    vl_logic;
        TDC_value_16    : out    vl_logic;
        TDC_value_15    : out    vl_logic;
        TDC_value_14    : out    vl_logic;
        TDC_value_13    : out    vl_logic;
        TDC_value_12    : out    vl_logic;
        TDC_value_11    : out    vl_logic;
        TDC_value_10    : out    vl_logic;
        TDC_value_9     : out    vl_logic;
        TDC_value_8     : out    vl_logic;
        TDC_value_7     : out    vl_logic;
        TDC_value_6     : out    vl_logic;
        TDC_value_5     : out    vl_logic;
        TDC_value_4     : out    vl_logic;
        TDC_value_3     : out    vl_logic;
        Q_31            : in     vl_logic;
        Q_30            : in     vl_logic;
        Q_29            : in     vl_logic;
        Q_28            : in     vl_logic;
        Q_27            : in     vl_logic;
        Q_26            : in     vl_logic;
        Q_25            : in     vl_logic;
        Q_24            : in     vl_logic;
        Q_23            : in     vl_logic;
        Q_22            : in     vl_logic;
        Q_21            : in     vl_logic;
        Q_20            : in     vl_logic;
        Q_19            : in     vl_logic;
        Q_18            : in     vl_logic;
        Q_17            : in     vl_logic;
        Q_16            : in     vl_logic;
        Q_15            : in     vl_logic;
        Q_14            : in     vl_logic;
        Q_13            : in     vl_logic;
        Q_12            : in     vl_logic;
        Q_11            : in     vl_logic;
        Q_10            : in     vl_logic;
        Q_9             : in     vl_logic;
        Q_8             : in     vl_logic;
        Q_7             : in     vl_logic;
        Q_6             : in     vl_logic;
        Q_5             : in     vl_logic;
        Q_4             : in     vl_logic;
        Q_3             : in     vl_logic;
        Q_2             : in     vl_logic;
        Q_1             : in     vl_logic;
        Q_110           : in     vl_logic;
        Q_210           : in     vl_logic;
        Q_32            : in     vl_logic;
        Q_41            : in     vl_logic;
        Q_51            : in     vl_logic;
        Q_61            : in     vl_logic;
        Q_71            : in     vl_logic;
        Q_81            : in     vl_logic;
        Q_91            : in     vl_logic;
        Q_101           : in     vl_logic;
        Q_111           : in     vl_logic;
        Q_121           : in     vl_logic;
        Q_131           : in     vl_logic;
        Q_141           : in     vl_logic;
        Q_151           : in     vl_logic;
        Q_161           : in     vl_logic;
        Q_171           : in     vl_logic;
        Q_181           : in     vl_logic;
        Q_191           : in     vl_logic;
        Q_201           : in     vl_logic;
        Q_211           : in     vl_logic;
        Q_221           : in     vl_logic;
        Q_231           : in     vl_logic;
        Q_241           : in     vl_logic;
        Q_251           : in     vl_logic;
        Q_261           : in     vl_logic;
        Q_271           : in     vl_logic;
        Q_281           : in     vl_logic;
        Q_291           : in     vl_logic;
        Q_301           : in     vl_logic;
        Q_311           : in     vl_logic;
        Q_112           : in     vl_logic;
        Q_212           : in     vl_logic;
        Q_33            : in     vl_logic;
        Q_42            : in     vl_logic;
        Q_52            : in     vl_logic;
        Q_62            : in     vl_logic;
        Q_72            : in     vl_logic;
        Q_82            : in     vl_logic;
        Q_92            : in     vl_logic;
        Q_102           : in     vl_logic;
        Q_113           : in     vl_logic;
        Q_122           : in     vl_logic;
        Q_132           : in     vl_logic;
        Q_142           : in     vl_logic;
        Q_152           : in     vl_logic;
        Q_162           : in     vl_logic;
        Q_172           : in     vl_logic;
        Q_182           : in     vl_logic;
        Q_192           : in     vl_logic;
        Q_202           : in     vl_logic;
        Q_213           : in     vl_logic;
        Q_222           : in     vl_logic;
        Q_232           : in     vl_logic;
        Q_242           : in     vl_logic;
        Q_252           : in     vl_logic;
        Q_262           : in     vl_logic;
        Q_272           : in     vl_logic;
        Q_282           : in     vl_logic;
        Q_292           : in     vl_logic;
        Q_302           : in     vl_logic;
        Q_312           : in     vl_logic;
        TDC_value_2     : out    vl_logic;
        TDC_value_1     : out    vl_logic;
        TDC_value_0     : out    vl_logic;
        Q_0             : in     vl_logic;
        Q_01            : in     vl_logic;
        Q_02            : in     vl_logic;
        enable_tdc      : in     vl_logic;
        devpor          : in     vl_logic;
        devclrn         : in     vl_logic;
        devoe           : in     vl_logic
    );
end TDC_result;
