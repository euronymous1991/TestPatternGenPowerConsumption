library verilog;
use verilog.vl_types.all;
entity Counter is
    port(
        Q_1             : out    vl_logic;
        Q_2             : out    vl_logic;
        Q_3             : out    vl_logic;
        Q_4             : out    vl_logic;
        Q_5             : out    vl_logic;
        Q_6             : out    vl_logic;
        Q_7             : out    vl_logic;
        Q_8             : out    vl_logic;
        Q_9             : out    vl_logic;
        Q_10            : out    vl_logic;
        Q_11            : out    vl_logic;
        Q_12            : out    vl_logic;
        Q_13            : out    vl_logic;
        Q_14            : out    vl_logic;
        Q_15            : out    vl_logic;
        Q_16            : out    vl_logic;
        Q_17            : out    vl_logic;
        Q_18            : out    vl_logic;
        Q_19            : out    vl_logic;
        Q_20            : out    vl_logic;
        Q_21            : out    vl_logic;
        Q_22            : out    vl_logic;
        Q_23            : out    vl_logic;
        Q_24            : out    vl_logic;
        Q_25            : out    vl_logic;
        Q_26            : out    vl_logic;
        Q_27            : out    vl_logic;
        Q_28            : out    vl_logic;
        Q_29            : out    vl_logic;
        Q_30            : out    vl_logic;
        Q_31            : out    vl_logic;
        OW1             : out    vl_logic;
        inst11          : in     vl_logic;
        system_reset    : in     vl_logic;
        inst10          : in     vl_logic;
        Q_0             : out    vl_logic;
        CLOCK_50        : in     vl_logic;
        devpor          : in     vl_logic;
        devclrn         : in     vl_logic;
        devoe           : in     vl_logic
    );
end Counter;
